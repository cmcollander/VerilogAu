// www.referencedesigner.com 
// Verilog Tutorial
// Hex to 7 Segment Example
 
module HexToInverseSevenSeg(
    input  [3:0]x,
    output reg [6:0]z
    );
    
    always @*
        case (x)
            4'b0000 : z = 7'b0000001;
            4'b0001 : z = 7'b1001111;
            4'b0010 : z = 7'b0010010; 
            4'b0011 : z = 7'b0000110;
            4'b0100 : z = 7'b1001100;
            4'b0101 : z = 7'b0100100;  
            4'b0110 : z = 7'b0100000;
            4'b0111 : z = 7'b0001111;
            4'b1000 : z = 7'b0000000;
            4'b1001 : z = 7'b0000100;
            4'b1010 : z = 7'b0001000; 
            4'b1011 : z = 7'b1100000;
            4'b1100 : z = 7'b0110001;
            4'b1101 : z = 7'b1000010;
            4'b1110 : z = 7'b0110000;
            4'b1111 : z = 7'b0111000;
        endcase
endmodule